//mux:4 to 1
`include "define.v"

module mux4(
    //input          clk,
    input   [31:0] pc_add4,
    input   [31:0] NOOP,
    input   [31:0] branch,
    input   [31:0] pc_jump,
    input   [1:0]  sel,
    output  reg [31:0] result
);
    initial begin
        result = 0;
    end
    always @(*) begin
        case (sel)
            `NextIns: result = pc_add4;
            `Jump: result = pc_jump;
            `Branch: result = branch;
            `NOOP: result = NOOP;
            default: result = pc_add4;
        endcase
    end
endmodule